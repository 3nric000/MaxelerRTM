XlxV61EB    1749     560a�e��Ҡx-���.�v�}܋R��� 	��{����F�n�A�j�@QuEߡ�VCR#h�ߎo~�S���L~�9&�
5��T�[p��ƟN�!��M�=Z������=2��4(��U�6�pRn��Tt��a���Q7AXe�}�&�|��C����)c��^�����ρT(V�.��˰B�m�]�P���w%��
P��%t��{/4O�J L>��n��_L�*T��#�Iu���eR�nÚ�G�@�f���X����G���9�z1K�z֟�&?���bHN��[!�ڸ)�5��cɍ{r�L���6����E��Y���bz���c;��Vj-p]�ۑi�{5V��q���������ڌ3q���#PrEã�Gf�'\���_p��/Onј�)���sN{��C�k��s:��7Մ����<C�:<ͺ���Sr�����fx��5���k0Sa+�ĉ��C�5��@��1{� gIo��@�����6��&��,��n!Te)�!Q�	�	�b�b"�h�?ix�!#n�%/��m�ַyA�`�*�^�<��ޜ`8^��Cb�%��|c�u
�!�m���킭�&����CJЂt��w�bn��)(�Q�;Q� �d�c�t9�.�HqFVLG2��ʯz�SD6�(��K��|��rb�cT����O�)�m�d�-	�O���3=e���.�4���A���ZF�6A�^9eP����΋̡���|^|낐�Y�vM��4�:�UQ_��4�"ʽ6d)��,�˱5�nGAI��fa"ױ�6T�������^ar��1�������ޝ��o��&�r@5=k��0@6���%��U����ė7�U�·����Y/S���E���v5T�7�f�[�vh(�
������]� WK�+�h!K;L�0��WG�(�I�o0.�>$�$���4h��91J�'�6lS��K�+&z��v'!�1eX|kfG��\Yz���%��[48�r�����s�,K�X���ѣ%�oQ�c6�9JU��c��6I�eF������R�83��	����gP ga�X��U�gBP�4����y~���aM�eU�K�LiVa�\7��bA��w�����
�GC�������Dr��@QF ��W�lN��AZ�5Q�rt�=�.�ݦ�L��I�q�9S��W-
oSbi���ZnM�Z�"�lc~H�|w��l` ��g'�%�7uF_컲�V�M�s�q�Ό��S�޹W�&Á����O��t6���ف��7����Z4x�����~��A'���u^R�$���o5��G�6�����Ŵ$��x�h�xm?�]M穓�qWj�f(l)N�?#��pc��4��w6#C����ΠD