XlxV61EB     3f3     1c06R6=��kKg��p������,�ͩ8�s���tOڣ|��(KR�T�I�Ɋ�^n��E�+r�v����D$��\���ī�J�%dKbd3��w4��  �*��:�5Fe�#t9���VU\bbb˦ѲoT�3���v�-���v��MY�?���7[~���Ől�nH:���p�U�pA�q��(�J�^$i����e5w�\�v�����^ӳq|�@E��7�kq5��+Q<��~ujsЯmޢ�Bb�+]��P|A��!(�[�u��63Ƽ�,�ѷf�T"Ē��~M嚷�aI�/��/�
���؎l�W��g-�h�ub�L�y�G�δsJ�GsN���H7B8rU`�i-wpl�!�!}�ua�x�y�»���I ���1��k����8d����]��f3#c��]�e���W�}�ۮ�eO��ӌ��