XlxV61EB    1623     670_^���
�9�\�NK2�U��_�����K�!��֣�f!�ݼ|����M`~-u��%P3nf<o�d���%u�ҾpM�n��"���7T�~�[�Q�K����۩|{���9t�H�nx�D�
��r+���׽��L����=���f��q�{|�IE�p�m:Ĵ�J*��lB�+<��/.�5�ֆك�l��.=:�2����T"ۅm1ٝ`��V�e���F�=�
zM���o�r�4�)<��S�����3��#C�IG	��
�XP�\`�J�;�n��-I��L̿R���$��B +5g��
f�7��3Ɖ0���ӷI�*�ʗ�f�M�sk� �X\���x���^��m0�]T�נ^��xC���[AZ!q9.���i�е�����tk��Wk{>�=G��ӮK����&�\��{�wf\�h����V�.�nk����Y���+���3��z<� �Z��B�ىb���͏�ݝ쿁#�⎭<^W�s���>*�N�`��o�No(�.���B�Ǻ{�遻�~����؟o+��]�}���3sҒ��W��Ɔ��N}p� ���yl���Y�h��d\>��0M%m�����u���7�Q����%�T�Q�,r�T��ʟ�7�V￝ߪN R5�AʜnB�p�1�{����@�4s�9���j�!�@��+��_-����#z���]*"op�	w�<�鳰�i��$���������~��VmRQ.�A�4� �j�\}�u������{r �������m9;�Hf��j���)���Vz��n3���1���_C$���nX�׏?�H�hTV�i�> ����T���_H!G~����9��93�L�IQ�5o��1H�('����'HZ+�7�#�t)@�m��7�W� �&��7!��2�U80��1�������4��@x҉�X��.]"��h���:$Bw�u5�pm���s��GO5?`{N�)����ڶ/�� ۴z ��cn��w��%.<��ΊhlL�����t�%y��qr�9�@�'�k˄�'X�_�'O��k,~��S�8aXTM�_����W�"Ј����f����=��X2�CD�n�6J>�\z���X�U��U�˓V��ޕ��oVk�0��M0Ƕ�t �q�Ig�'�AU^�BA�ߤط]υt��Iobʇ�Z�H�A�N����Y� <�a0�GB(�T��@������+q�C��/�үJ?E�7������X��r@�i��6F�hC���7n�õ��$j���<_�-7ͱ`�$�D�|-" /�?bC����B���X����58�])n�!Z/����q.��k����^-����c�f�(gS3�O�y30\�ͣ�IG��ƶ�v�yrݚ��ۏ��b��Q��W��ܠ���O_�S�R�l��Lե����S�`
�*_\�f�H��!Nsi���q�|�2V�����O��ɍr� �7�^���wd�p���:@�2�0=9�Q��ƌuB���ID$u7ڮ
s��蟓գƩ�C&�>�!@�����`�� ��
tP4$U�:&�U�OS���A�֥ȍLS�Vdy_
�Ƴ�0z�B���5^�U����,��$�lVD�
��+��� �T
K�%Y�4Q�륎��\q���@�ZEl�XC2�