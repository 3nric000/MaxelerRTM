XlxV61EB     9c1     2e0�pb�T�����WW��-���ƤƢ��pE�;����3d�^�R�8d�ǆǘ}˪�4�i�s|�2A�����=�.�g����  �|�{;��<�Q�399��78���qH'����1>���8�Hl�������$F/C}�$"�ȉlI��ȋt�M�L����AN��Gx�N�����"��$=� ua=
Չ���w~�:����+��d�i6�ȵ>h�ٖA�sNbI�I��6���d�ϵ ��hHr�$���M7���	������0������r�PVz;G���n��Y~AT1��c�6��\����,��.ru��Vn ���8d�%���+�}�0�.t)��䦸;���(B�I�$��Sy�/� �Q����$ýE��P0�_�k�`wʌ�k���,�b̡{��r���5�:x��;��[YL�e4$I+@4=Eӑ�b�~Z�Z?�n�#q��[�_z2s(r`�.��s�1�L�uOJ�Q(�j��y��X���vz�Q$�<��0��DG�h�jJu�ھ~

yל!w�ւ(�<Q}|�v(m���}�w�6�;W� U�=��� �J����O�{`���5�}�����4z]�_��
 &|u��^C����� 6V���)hf�1H45�1�]o��HT��lMjv"2�g�V��kJ?���k�;�gƒ�˚��-�pT��7����1AH3}a�)���  ���?�bZ	�