XlxV61EB    2aeb     790� �����3�b
hֶ���gM�c	J�<���N{H��jdjn��7�m�ui���W/�]�^�%`1����ķ���MP쬅E�Ƹ�9�R�&�$ƕsR7��C�_���������rm�>��� OQ/��S$]�"���m���e϶�唙t�y���<{lp"�	�L�8
��vi�0:�τZb|Q����4�J�Q�+��Ec�~7�L� ɘ/�a�YTD�ZD}d��}W�)���E����T`���N0W�����'�y���ީ�-s�̵n���P��	�O!�Tkt2v���>�˻�t��K���2S���_&���rH|`�� �g����L��\o7�w�o�x�W��x 8��Df�t8G�2ΜQbn<��N�֗h�r���_k7mR�lJ̈́����"��h�0Pr��܁�MĞ�K���-It+w�7�7��-#���D�*[�c�<F��x龈��������w8D���������iU�EjK�F�!ܦҍ�0���1�_�vr�T��4�P��e3�ai^&�W5*@��\fUqST� �	<��ۮ����"섆G��A)�W�����/i����}�Vnu�@-of0�v˶^���2�Q�Vv���ߢѪ�B�w/�X3�-�血`�5EgZ��bA;g����u@���o�;�$�o� 0���9�'��CT�-�ص�q�
�����j��*{"�������R�J'u�YLq$�ѳ��j��3�F!��Wf$��^	m��ᐮ��̗&��4F�Ã�e���J��<���B�H�i���~��Ȩ���Ӳ0e���m�}��C��������<d�+�1|����7�?��,.#?�TJ:�3�I��'wrL#��^�O(�f�7�C�?tD��E,~�c��`d��Yl���;`�9�4HƄ��+�&��~�Qr�47x�ٴƝK|�.����Sn')�����Ί��A��˷���TԔ�T^���ϫ'�'SH4��R�q�$c$���)���:���^��R�tnw1��8��M��1�'t�30�q����e�oE�:G�J��#NJ��a�X��V	�4}AɢY8�"�S-�̺^o�1��!d��J;4)V,D��?bA�����И�N'�Uˈ��^KL�p������J�� +g��'Ʀ��I+��<���Vv��ZZl65r��	.�f���{��̘h-�R��{�WsĽ-�_c���=��K�D9���m�b���q��m5پn�L�iu}� ���>� ��tܮQ����L�M���mȘ�yc��d\f�X2|g=��u���&u��\Ι�0�=솈��-���A��PU�n\�o��S���~��
A��&h�Ly��{�b��"721��A_^����O���i�"}>��}G�M%�hpJJ.r����\�}��Eٔ�(��G��i�����%MgWY=3h&Dzj,XzY=uS)J�%����q�wE �p$@�yc�M�!��k��K��۲܌@s�G_��(��b���|��-��a �8�#�э���~P�
Pn5�M-��ƕ3��,��9%�@��
u`��#"M�@ۈ%��dt��#�� �oEd��Ta�{�[P�d�n=p�Ai$\����n	W^���_f�,"�E���WWNX?�#CW�sv˨K�����!�$���<���J�KcA�.��&1LD�$W�(&�B��?����4��:Е��z���.d��Oa�w�Ø�
�$�xi�C����yw��5w���'�Q=6�\��R9�\9������ģY����4��w[��#{"�)K��H��rn�Tq_[qs���f�J?@�l (�Z�TK�e�p���=�|w����uÙTR/
<�s=4hr���.�$ A
R54HTJ� GS�!q�)�&q��:<�_E
�|�S��