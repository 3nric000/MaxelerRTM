XlxV61EB    1c81     7e0�LG3����y49��8��41n�q�G��H,�8�5��iu=��M��U
Yǜ,��?=�ʄh@��?'�;3Z9 �E{��,sN�vnM-,����M.4 5�s��I��C��'�h+vCM&&�u��S�]���r��v��ۭ��L�=��5!u�܋]� �ˀ�� I# ",�ӕ�UQ������7Q����w(�{��EKf�m%O�Zy:���ܓ)攀JUW�2���gA�|��Ee��G`gZ|s�3�\�~��\�v��5:�����vL�id��#�Qd�K]���09B��G*��*G��>�sA��T˄���	�'@SHX���A,���N��So�>&؍<�32�W��rR�4��|F���lf���,%��2Q�*<��k�ť�ABFP~��ixiqcb (;Z��M7m�d��J�?�e�>����0I�Ώ��,wP7�<��yw�,�)T�0�J��A�F��"�ͽM���l�E}R�^Ee�`�}�V���F�����A�α����3�7��.���ɽκ��J�����{�e�Y�!�q�v��6�^Xp�k�F<0"�I�_&�Qp���G��4G�V����Jk�`��q��0*���meɕt��D}ÄI ���v���ay�|��R�#D�3�2u�i����Ҷ����V���4���8ғ�ki�l'���ti���$��i�'����!��7�ЋcI�Ŕ��<��\-T=�Zj	�	cy��O��k˄]h��?��h��e =X`�W0X�0P��-�e*����y*k�<=;���C���J�����Ug��cȋ������''�-Y�ŏ]�oиR�P���DI�:R���Ж���	�fH����<y�����pj��$��;�2�z�X&�¾=��S���J��I��0Ǣg�4�|��	��_Jc��`��qKU�s\eU��Յ�����*�#�!��g�%��N@XU�α��y��@+�s�Fh<OU����0yV����د��3ϵ]_�JC�&)���D@?�*{��G����z�n\��iZ_��J.\�L{��/V+��q�u�ԭ���|�^�L�h�z_j:�NV�Ց޳�ԥ��d��W�,���6Zg9�m'����E��%�&����v{�nC��_�N���馪�Wd׀��E�����
d}�������4��R����3ٚoHe:��M�>��&�/kb��r���� ��6s�q��e������S3"���o������FrS�ي�%oV��b�~p\���ll��KH����<�$�љA�(���u��s����lc�F֒�y�-Ɣ'��v�q��	�q�è��\N����_�홵�EC$d���dS�z�����"�e���sr����`&�"�P=�E'ݮ���"�k��[��������a�]���x1X�ܝ3sXj�D���uDek�ɇKv��zhh�ؤ/�ߨ�-��� �OW6�&}�B�+��X:���lHK��Ţβ�?�6�6Q/M�����ػ����V�w�����o3��S0yk�h����B�m(�T|^ذ1��Qĸ�ܛN1��F�,uS��n)�'��g����:GQ��)Cd�dc�I{s�
�3z�bi�2����7 N8Úze��LU(�if35k	������-�M������|��/���t�q�,3yUij+��q�r�H��4�t!��
M>�J'�FH-��o�b(%�ȯ�j��r~{��{6z�v�C� ]���62A�s5��ݰ���T�C�{n��?FWT��V��VFG��C�������Ҹڈ���$������=^��� ���t�7�#w	J�H�<:^ �ڜ9Ȍ��$,]��+hCyN I/4�M���q6>8������\����םfBs �s��نts�W�S�v�� ��lL���3q1�z���9��Y����b�c(_�׻�K͢�fW}��S�8 ��v 